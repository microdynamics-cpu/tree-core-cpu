module hello;
   initial begin 
      $display("Hello World");
      $finish; 
   end
endmodule
